`timescale 1ns / 1ps

module logic_func0_tb;

    reg  A, B, C, D;
    wire F0;

    integer errors;
    integer i;
    reg expected;

    // Instantiate the Unit Under Test (UUT)
    logic_func0 uut (
        .p(A),
        .q(B),
        .r(C),
        .s(D),
        .F0(F0)
    );

    initial begin
        errors = 0;

        $display("===========================================");
        $display("   Logic Func0 Testbench - Starting Tests");
        $display("===========================================");
        $display("   Testing: F0 = (A & B) | (C & D)");
        $display("===========================================");

        for (i = 0; i < 16; i = i + 1) begin
            {A, B, C, D} = i[3:0];
            #10;
            expected = (A & B) | (C & D);
            if (F0 !== expected) begin
                $display("FAIL: A=%b, B=%b, C=%b, D=%b, F0=%b (expected %b)", A, B, C, D, F0, expected);
                errors = errors + 1;
            end else begin
                $display("PASS: A=%b, B=%b, C=%b, D=%b, F0=%b", A, B, C, D, F0);
            end
        end

        $display("===========================================");
        if (errors == 0) begin
            $display("   ALL TESTS PASSED!");
            $display("===========================================");
            $finish;
        end else begin
            $display("   TESTS FAILED: %0d errors", errors);
            $display("===========================================");
            $fatal(1, "Testbench failed");
        end
    end

endmodule
